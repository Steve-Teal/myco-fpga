---------------------------------------------------------------------
--
-- Built with PASM version 1.3
-- File name: myco_mem.vhd
-- 6-12-2020 18:54:47
-- 
---------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity myco_mem is
port (
    clock        : in std_logic;
    clock_enable : in std_logic;
    address      : in std_logic_vector(9 downto 0);
    data_out     : out std_logic_vector(15 downto 0);
    data_in      : in std_logic_vector(15 downto 0);
    write_enable : in std_logic);
end entity;

architecture rtl of myco_mem is

    type ram_type is array (0 to 1023) of std_logic_vector(15 downto 0);
    signal ram : ram_type := (
			X"B012",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0001",X"0002",
			X"0003",X"0004",X"0222",X"1001",X"1002",X"1003",X"1004",X"1006",
			X"1007",X"A011",X"A00E",X"900D",X"100C",X"5223",X"D029",X"1005",
			X"A00E",X"0224",X"A010",X"E0A5",X"E041",X"E04F",X"0005",X"2225",
			X"B01F",X"0222",X"1005",X"E0A5",X"0226",X"2009",X"4227",X"1030",
			X"B031",X"B0AF",X"B0B2",X"B0B5",X"B0CB",X"B0CE",X"B0D1",X"B105",
			X"B131",X"B17E",X"B183",X"B186",X"B18B",X"B190",X"B1DC",X"B1DF",
			X"B0AF",X"0009",X"A00E",X"E082",X"D04E",X"0222",X"1009",X"A00E",
			X"E05D",X"E082",X"D04E",X"0009",X"2225",X"B046",X"F000",X"0008",
			X"A00E",X"E082",X"D05C",X"0222",X"1008",X"A00E",X"E05D",X"E082",
			X"D05C",X"0008",X"2225",X"B054",X"F000",X"0009",X"100B",X"E086",
			X"4008",X"100A",X"E07C",X"000A",X"100B",X"E075",X"7005",X"0228",
			X"C06A",X"0229",X"500A",X"400B",X"100A",X"7005",X"522A",X"222B",
			X"422C",X"1073",X"000A",X"B074",X"F000",X"7005",X"522A",X"222B",
			X"1079",X"B07A",X"100A",X"F000",X"7005",X"C07F",X"F000",X"800A",
			X"100A",X"F000",X"E093",X"3225",X"C082",X"F000",X"E089",X"E089",
			X"E089",X"000B",X"200B",X"100B",X"F000",X"E090",X"E090",X"E090",
			X"700A",X"100A",X"F000",X"900D",X"600C",X"D098",X"0222",X"F000",
			X"100A",X"022D",X"A010",X"900D",X"600C",X"600A",X"D096",X"000A",
			X"600C",X"100C",X"622E",X"500A",X"F000",X"E075",X"E07C",X"000A",
			X"522F",X"1008",X"E08D",X"000A",X"522F",X"1009",X"F000",X"0005",
			X"2225",X"B02A",X"0008",X"A00E",X"B0AF",X"0230",X"2008",X"10B8",
			X"B0B9",X"A010",X"B0AF",X"0001",X"0002",X"0005",X"000A",X"0014",
			X"0032",X"0064",X"00C8",X"01F4",X"03E8",X"07D0",X"1388",X"2710",
			X"4E20",X"7530",X"EA60",X"0005",X"3008",X"B02A",X"0008",X"1001",
			X"B0AF",X"0231",X"2008",X"4227",X"10D6",X"0001",X"B0D7",X"B0AF",
			X"B0E8",X"B0EA",X"B0EC",X"B0EE",X"B0F0",X"B0F2",X"B0F4",X"B0F6",
			X"B103",X"B0AF",X"B0AF",X"B0AF",X"B0AF",X"B0AF",X"B0AF",X"B0AF",
			X"1002",X"B0AF",X"1003",X"B0AF",X"1004",X"B0AF",X"A00E",X"B0AF",
			X"0225",X"B0F7",X"0223",X"B0F7",X"0232",X"B0F7",X"0233",X"100A",
			X"7001",X"C0FD",X"900E",X"400A",X"B0EE",X"000A",X"622F",X"100A",
			X"900E",X"500A",X"B0EE",X"A011",X"B0AF",X"0234",X"2008",X"4227",
			X"110A",X"900F",X"B10B",X"B0AF",X"B11B",X"B11E",X"B120",X"B122",
			X"B124",X"B126",X"B128",X"B12A",X"B12F",X"B12F",X"B0AF",X"B0AF",
			X"B0AF",X"B0AF",X"B0AF",X"0002",X"1001",X"B0AF",X"0003",X"B11C",
			X"0004",X"B11C",X"900F",X"B11C",X"5225",X"B12B",X"5223",X"B12B",
			X"5232",X"B12B",X"5233",X"D12D",X"B11C",X"0225",X"B11C",X"0222",
			X"B11C",X"0235",X"2008",X"4227",X"1136",X"0001",X"B137",X"B0AF",
			X"B147",X"B14A",X"B14C",X"B14E",X"B150",X"B164",X"B176",X"B178",
			X"B17A",X"B17C",X"B0AF",X"B0AF",X"B0AF",X"B0AF",X"B0AF",X"2225",
			X"1001",X"B0AF",X"3225",X"B148",X"2002",X"B148",X"3002",X"B148",
			X"0002",X"100B",X"E086",X"0232",X"100A",X"000B",X"200B",X"100B",
			X"5236",X"D15B",X"B15E",X"000B",X"2001",X"100B",X"000A",X"3225",
			X"D154",X"000B",X"522F",X"B148",X"0002",X"100B",X"E086",X"0232",
			X"100A",X"0001",X"2001",X"1001",X"300B",X"C170",X"4225",X"1001",
			X"000A",X"3225",X"D168",X"0001",X"522F",X"B148",X"5002",X"B148",
			X"4002",X"B148",X"6002",X"B148",X"622F",X"B148",X"0008",X"100B",
			X"E086",X"1006",X"B0AF",X"0006",X"4008",X"B02A",X"0003",X"3225",
			X"C0AF",X"1003",X"B183",X"0004",X"3225",X"C0AF",X"1004",X"B183",
			X"0237",X"2008",X"4227",X"1194",X"B195",X"B0AF",X"B1A5",X"B1A9",
			X"B1AD",X"B1B1",X"B1B3",X"B1B5",X"B1B7",X"B1BD",X"B1BF",X"B1C1",
			X"B1C3",X"B1C9",X"B1CD",X"B1D1",X"B1D5",X"0002",X"3001",X"C1D9",
			X"B0AF",X"0001",X"3002",X"C1D9",X"B0AF",X"0001",X"3002",X"D0AF",
			X"B1D9",X"0225",X"B1B8",X"0223",X"B1B8",X"0232",X"B1B8",X"0233",
			X"100B",X"900F",X"500B",X"D1D9",X"B0AF",X"0225",X"B1C4",X"0223",
			X"B1C4",X"0232",X"B1C4",X"0233",X"100B",X"900F",X"500B",X"D0AF",
			X"B1D9",X"900D",X"5225",X"D0AF",X"B1D9",X"900D",X"5223",X"D0AF",
			X"B1D9",X"900D",X"5225",X"D1D9",X"B0AF",X"900D",X"5223",X"D1D9",
			X"B0AF",X"0005",X"2223",X"B02A",X"0005",X"1007",X"B183",X"0007",
			X"1005",X"B0AF",X"6451",X"4E80",X"C398",X"8295",X"4D80",X"C39E",
			X"829A",X"4B81",X"C394",X"8390",X"4781",X"C39A",X"8394",X"4382",
			X"C390",X"8490",X"1128",X"1828",X"3471",X"5459",X"2634",X"6954",
			X"5926",X"34FF",X"54CE",X"7133",X"22CC",X"3240",X"2271",X"54CE",
			X"3439",X"FFFF",X"86D0",X"4071",X"5423",X"CD34",X"D840",X"543B",
			X"FFFF",X"FFFF",X"4F93",X"4553",X"1911",X"2119",X"1121",X"1911",
			X"20B4",X"10E0",X"23CE",X"3223",X"CC31",X"E0FF",X"23CF",X"3223",
			X"CD31",X"E0FF",X"CC31",X"4054",X"23CE",X"32CF",X"E0CC",X"3371",
			X"23CC",X"313C",X"0000",X"0002",X"012C",X"0001",X"0031",X"B000",
			X"00FF",X"FF00",X"003F",X"01E2",X"1000",X"001E",X"0003",X"000F",
			X"00BB",X"00D7",X"0004",X"0008",X"010B",X"0137",X"0100",X"0195",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
			X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000");
begin

    process(clock)
    begin
        if rising_edge(clock) then
            if clock_enable = '1' then
                if write_enable = '1' then
                    ram(to_integer(unsigned(address))) <= data_in;
                else
                    data_out <= ram(to_integer(unsigned(address)));
                end if;
            end if;
        end if;
    end process;

end rtl;

--- End of file ---
